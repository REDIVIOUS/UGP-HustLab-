//verilint 143 sticky_off
`define NUM_CORES 1
`define MIPS_CMP_NUM_CORES 1
`define MIPS_CORE0_MODULE core
`define MIPS_CORE0_PRESENT 1
`define MIPS_UNIQUIFIDE_CORE_SYSTEM 0
`define MIPS_CMP_MODULE mips_cmp_stub
`define MIPS_L2_MODULE mips_l2_stub
`define MIPS_SC_MODULE mips_sc_stub
`define MIPS_PROJECT_M14KEc 1
//verilint 143 on
